library ieee;
use ieee.std_logic_1164.all;

package tb_pkg is

  signal clk : std_logic := '0';

end package tb_pkg;
